// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Author: Florian Zaruba, ETH Zurich
// Date: 19.03.2017
// Description: Test-harness for Ariane
//              Instantiates an AXI-Bus and memories

`include "axi/assign.svh"
`include "register_interface/typedef.svh"
`include "register_interface/assign.svh"
`define PMU_BLOCK

module cva6_subsystem 
  import axi_pkg::xbar_cfg_t;
  import ariane_soc::*;
  import udma_subsystem_pkg::N_CAN;  
#(
  parameter int unsigned AXI_USER_WIDTH    = 1,
  parameter int unsigned AXI_ADDRESS_WIDTH = 64,
  parameter int unsigned AXI_DATA_WIDTH    = 64,
`ifdef PMU_BLOCK
  parameter int unsigned PMU_NUM_COUNTER   = 64,
`endif
`ifdef DROMAJO
  parameter bit          InclSimDTM        = 1'b0,
`else
  parameter bit          InclSimDTM        = 1'b1,
`endif
  parameter int unsigned NUM_WORDS         = 2**25,         // memory size
  parameter bit          StallRandomOutput = 1'b0,
  parameter bit          StallRandomInput  = 1'b0,
  parameter bit          JtagEnable        = 1'b1
) (
  input  logic             clk_i,
  input  logic             rtc_i,
  input  logic             rst_ni,
  input  logic             sync_rst_ni,
  input  logic             cva6_clk_i,
  input  logic             cva6_rst_ni,
  output logic             dm_rst_o,
  input  logic [31*4-1:0]  udma_events_i,
  input  logic             c2h_irq_i,
  input  logic             cluster_eoc_i,
  input  logic [N_CAN-1:0] can_irq_i,
  input  logic             cl_dma_pe_evt_i,
  input  logic             dmi_req_valid,
  output logic             dmi_req_ready,
  input  logic [ 6:0]      dmi_req_bits_addr,
  input  logic [ 1:0]      dmi_req_bits_op,
  input  logic [31:0]      dmi_req_bits_data,
  output logic             dmi_resp_valid,
  input  logic             dmi_resp_ready,
  output logic [ 1:0]      dmi_resp_bits_resp,
  output logic [31:0]      dmi_resp_bits_data,
  // JTAG
  input  logic             jtag_TCK,
  input  logic             jtag_TMS,
  input  logic             jtag_TDI,
  input  logic             jtag_TRSTn,
  output logic             jtag_TDO_data,
  output logic             jtag_TDO_driven,

  `ifdef PMU_BLOCK
  output pmu_pkg::pmu_event_t spu_core_0_out,
  output pmu_pkg::pmu_event_t spu_core_1_out,
  output pmu_pkg::pmu_event_t spu_core_2_out,
  output pmu_pkg::pmu_event_t spu_core_3_out,
  // From AXI4-Lite Bar
  AXI_BUS.Slave               axi_lite_slave,
  // PMU Interrupt Signal
  input  logic [PMU_NUM_COUNTER-1:0]  pmu_intr_i,
  `endif

  //SERIAL LINK
  output ser_link_to_pad serial_link_to_pad,
  input  pad_to_ser_link pad_to_serial_link,
  REG_BUS.in             serial_linkcfg_reg_master,

  // CVA6 DEBUG UART
  input  logic            cva6_uart_rx_i,
  output logic            cva6_uart_tx_o,

  AXI_BUS.Master          axi_lite_master,
  AXI_BUS.Master          l2_axi_master,
  AXI_BUS.Master          apb_axi_master,
  AXI_BUS.Master          hyper_axi_master,
  AXI_BUS.Master          cluster_axi_master,
  AXI_BUS.Slave           cluster_axi_slave
);
     // disable test-enable
  logic        test_en;
  logic        ndmreset;
  logic        ndmreset_n;
  logic [3:0]       debug_req_core;
  
  logic        jtag_enable;
  logic        init_done;

  logic        debug_req_valid;
  logic        debug_req_ready;
  logic        debug_resp_valid;
  logic        debug_resp_ready;

  logic        jtag_req_valid;
  logic [6:0]  jtag_req_bits_addr;
  logic [1:0]  jtag_req_bits_op;
  logic [31:0] jtag_req_bits_data;
  logic        jtag_resp_ready;
  logic        jtag_resp_valid;

  dm::dmi_req_t  jtag_dmi_req;
  dm::dmi_req_t  dmi_req;

  dm::dmi_req_t  debug_req;
  dm::dmi_resp_t debug_resp;

  assign test_en = 1'b0;
  assign jtag_enable = JtagEnable;
   
  AXI_BUS_ASYNC_GRAY #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH   ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH      ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH      ),
    .LOG_DEPTH      ( 1                   )
  ) cva6_axi_master_dst_0();

  AXI_BUS_ASYNC_GRAY #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH   ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH      ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH      ),
    .LOG_DEPTH      ( 1                   )
  ) cva6_axi_master_dst_1();

  AXI_BUS_ASYNC_GRAY #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH   ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH      ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH      ),
    .LOG_DEPTH      ( 1                   )
  ) cva6_axi_master_dst_2();

  AXI_BUS_ASYNC_GRAY #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH   ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH      ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH      ),
    .LOG_DEPTH      ( 1                   )
  ) cva6_axi_master_dst_3();

  AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH   ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH      ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH      )
  ) slave[ariane_soc::NrSlaves-1:0]();

  AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH   ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH      ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH      )
  ) slave_to_spu[ariane_soc::NumCores-1:0]();
 
  AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH   ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH      ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH      )
  ) serial_link_master();

  AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH   ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH      ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH      )
  ) serial_link_cut();
   
  AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
  ) master[ariane_soc::NB_PERIPHERALS-1:0]();

  AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
  ) hyper_axi_master_cut();

  AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
  ) hyper_axi_master_redirect();

  AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
  ) cluster_axi_master_cut();
  
  assign ndmreset_n = sync_rst_ni;
   
  // ------------------------------
  // AXI4-Lite Master to AXI4 Slave
  // ------------------------------

  ariane_axi_soc::req_t   dummy_req;                                
  ariane_axi_soc::resp_t  dummy_resp;
  // assign dummy_req  = '0;
  // assign dummy_resp = '0;

  `ifdef PMU_BLOCK
    `AXI_ASSIGN ( slave[ariane_soc::AXI4_Lite], axi_lite_slave )
  `else
    `AXI_ASSIGN_FROM_REQ ( slave[ariane_soc::AXI4_Lite], dummy_req  )
    `AXI_ASSIGN_TO_RESP  ( dummy_resp, slave[ariane_soc::AXI4_Lite] )
  `endif 

  // ---------------
  // Debug
  // ---------------
  assign init_done = rst_ni;
   
  initial begin
    if (riscv::XLEN != 32 & riscv::XLEN != 64) $error("XLEN different from 32 and 64");
  end

  // debug if MUX
  assign debug_req_valid     = (jtag_enable) ? jtag_req_valid     : dmi_req_valid;
  assign debug_resp_ready    = (jtag_enable) ? jtag_resp_ready    : dmi_resp_ready;
  assign debug_req           = (jtag_enable) ? jtag_dmi_req       : dmi_req;
  assign jtag_resp_valid     = (jtag_enable) ? debug_resp_valid   : 1'b0;
  assign dmi_resp_valid      = (jtag_enable) ? 1'b0               : debug_resp_valid;

  dmi_jtag  #(
    .IdcodeValue ( 32'h20001001)
    ) i_dmi_jtag (
    .clk_i            ( clk_i           ),
    .rst_ni           ( rst_ni          ),
    .testmode_i       ( test_en         ),
    .dmi_req_o        ( jtag_dmi_req    ),
    .dmi_req_valid_o  ( jtag_req_valid  ),
    .dmi_req_ready_i  ( debug_req_ready ),
    .dmi_resp_i       ( debug_resp      ),
    .dmi_resp_ready_o ( jtag_resp_ready ),
    .dmi_resp_valid_i ( jtag_resp_valid ),
    .dmi_rst_no       (                 ), // not connected
    .tck_i            ( jtag_TCK        ),
    .tms_i            ( jtag_TMS        ),
    .trst_ni          ( jtag_TRSTn      ),
    .td_i             ( jtag_TDI        ),
    .td_o             ( jtag_TDO_data   ),
    .tdo_oe_o         ( jtag_TDO_driven )
  );

  assign dmi_req_ready = debug_req_ready ;    
  assign dmi_req.addr = dmi_req_bits_addr;
  assign dmi_req.data = dmi_req_bits_data;
  // SiFive's SimDTM Module
  // Converts to DPI calls
  assign dmi_req.op = dm::dtm_op_e'(dmi_req_bits_op);

  assign dmi_resp_bits_data = debug_resp.data;
  assign dmi_resp_bits_resp = debug_resp.resp;

  // this delay window allows the core to read and execute init code
  // from the bootrom before the first debug request can interrupt
  // core. this is needed in cases where an fsbl is involved that
  // expects a0 and a1 to be initialized with the hart id and a
  // pointer to the dev tree, respectively.
  localparam int unsigned DmiDelCycles = 500;

  logic [3:0] debug_req_core_ungtd;
  int dmi_del_cnt_d, dmi_del_cnt_q;

  assign dmi_del_cnt_d  = (dmi_del_cnt_q) ? dmi_del_cnt_q - 1 : 0;
  assign debug_req_core = (dmi_del_cnt_q) ? 1'b0 : debug_req_core_ungtd;

  always_ff @(posedge clk_i or negedge rst_ni) begin : p_dmi_del_cnt
    if(!rst_ni) begin
      dmi_del_cnt_q <= DmiDelCycles;
    end else begin
      dmi_del_cnt_q <= dmi_del_cnt_d;
    end
  end

  ariane_axi_soc::req_t    dm_axi_m_req;
  ariane_axi_soc::resp_t   dm_axi_m_resp;

  logic                dm_slave_req;
  logic                dm_slave_we;
  logic [64-1:0]       dm_slave_addr;
  logic [64/8-1:0]     dm_slave_be;
  logic [64-1:0]       dm_slave_wdata;
  logic [64-1:0]       dm_slave_rdata;

  logic                dm_master_req;
  logic [64-1:0]       dm_master_add;
  logic                dm_master_we;
  logic [64-1:0]       dm_master_wdata;
  logic [64/8-1:0]     dm_master_be;
  logic                dm_master_gnt;
  logic                dm_master_r_valid;
  logic [64-1:0]       dm_master_r_rdata;

  // debug module
  dm_top #(
    .NrHarts              ( 4                           ),
    .BusWidth             ( AXI_DATA_WIDTH              )
    // .SelectableHarts      ( 1'b1                        )
  ) i_dm_top (
    .clk_i                ( clk_i                       ),
    .rst_ni               ( rst_ni                      ), // PoR
    .testmode_i           ( test_en                     ),
    .ndmreset_o           ( dm_rst_o                    ),
    .dmactive_o           (                             ), // active debug session
    .debug_req_o          ( debug_req_core_ungtd        ),
    .unavailable_i        ( '0                          ),
    .hartinfo_i           ( {4{ariane_pkg::DebugHartInfo}} ),
    .slave_req_i          ( dm_slave_req                ),
    .slave_we_i           ( dm_slave_we                 ),
    .slave_addr_i         ( dm_slave_addr               ),
    .slave_be_i           ( dm_slave_be                 ),
    .slave_wdata_i        ( dm_slave_wdata              ),
    .slave_rdata_o        ( dm_slave_rdata              ),
    .master_req_o         ( dm_master_req               ),
    .master_add_o         ( dm_master_add               ),
    .master_we_o          ( dm_master_we                ),
    .master_wdata_o       ( dm_master_wdata             ),
    .master_be_o          ( dm_master_be                ),
    .master_gnt_i         ( dm_master_gnt               ),
    .master_r_valid_i     ( dm_master_r_valid           ),
    .master_r_rdata_i     ( dm_master_r_rdata           ),
    .dmi_rst_ni           ( rst_ni                      ),
    .dmi_req_valid_i      ( debug_req_valid             ),
    .dmi_req_ready_o      ( debug_req_ready             ),
    .dmi_req_i            ( debug_req                   ),
    .dmi_resp_valid_o     ( debug_resp_valid            ),
    .dmi_resp_ready_i     ( debug_resp_ready            ),
    .dmi_resp_o           ( debug_resp                  )
  );


  axi2mem #(
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
  ) i_dm_axi2mem (
    .clk_i      ( clk_i                     ),
    .rst_ni     ( rst_ni                    ),
    .slave      ( master[ariane_soc::Debug] ),
    .req_o      ( dm_slave_req              ),
    .we_o       ( dm_slave_we               ),
    .addr_o     ( dm_slave_addr             ),
    .be_o       ( dm_slave_be               ),
    .data_o     ( dm_slave_wdata            ),
    .data_i     ( dm_slave_rdata            )
  );

  `AXI_ASSIGN_FROM_REQ(slave[ariane_soc::DEBUG],dm_axi_m_req)
  `AXI_ASSIGN_TO_RESP(dm_axi_m_resp,slave[ariane_soc::DEBUG])


   
  axi_adapter #(
    .DATA_WIDTH            ( AXI_DATA_WIDTH            ),
    .AXI_ID_WIDTH          ( ariane_soc::IdWidth       )
  ) i_dm_axi_master (
    .clk_i                 ( clk_i                     ),
    .rst_ni                ( rst_ni                    ),
    .req_i                 ( dm_master_req             ),
    .type_i                ( ariane_axi::SINGLE_REQ    ),
    .busy_o                (                           ),
    .gnt_o                 ( dm_master_gnt             ),
    .gnt_id_o              (                           ),
    .addr_i                ( dm_master_add             ),
    .we_i                  ( dm_master_we              ),
    .wdata_i               ( dm_master_wdata           ),
    .be_i                  ( dm_master_be              ),
    .size_i                ( 2'b11                     ), // always do 64bit here and use byte enables to gate
    .id_i                  ( '0                        ),
    .valid_o               ( dm_master_r_valid         ),
    .rdata_o               ( dm_master_r_rdata         ),
    .id_o                  (                           ),
    .critical_word_o       (                           ),
    .critical_word_valid_o (                           ),
    .axi_req_o             ( dm_axi_m_req              ),
    .axi_resp_i            ( dm_axi_m_resp             )
  );


  // ---------------
  // ROM
  // ---------------
  logic                         rom_req;
  logic [AXI_ADDRESS_WIDTH-1:0] rom_addr;
  logic [AXI_DATA_WIDTH-1:0]    rom_rdata;

  axi2mem #(
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
  ) i_axi2rom (
    .clk_i  ( clk_i                   ),
    .rst_ni ( ndmreset_n              ),
    .slave  ( master[ariane_soc::ROM] ),
    .req_o  ( rom_req                 ),
    .we_o   (                         ),
    .addr_o ( rom_addr                ),
    .be_o   (                         ),
    .data_o (                         ),
    .data_i ( rom_rdata               )
  );

`ifdef DROMAJO
  dromajo_bootrom i_bootrom (
    .clk_i      ( clk_i     ),
    .req_i      ( rom_req   ),
    .addr_i     ( rom_addr  ),
    .rdata_o    ( rom_rdata )
  );
`else
  bootrom i_bootrom (
    .clk_i      ( clk_i     ),
    .req_i      ( rom_req   ),
 `ifdef FPGA_EMUL
    .rst        ( ndmreset_n),
 `endif                   
    .addr_i     ( rom_addr  ),
    .rdata_o    ( rom_rdata )
  );
`endif

  // ---------------
  // AXI L2 Slave
  // ---------------

  axi_riscv_atomics_wrap #(
    .AXI_ADDR_WIDTH     ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH     ( AXI_DATA_WIDTH           ),
    .AXI_ID_WIDTH       ( ariane_soc::IdWidthSlave ),
    .AXI_USER_WIDTH     ( AXI_USER_WIDTH           ),
    .AXI_MAX_READ_TXNS  ( 8                        ),
    .AXI_MAX_WRITE_TXNS ( 8                        ),
    .RISCV_WORD_WIDTH   ( 64                       )
  ) i_axi_riscv_atomicsl2 (
    .clk_i,
    .rst_ni ( ndmreset_n                ),
    .slv    ( master[ariane_soc::L2SPM] ),
    .mst    ( l2_axi_master             )
  );

  // ---------------
  // AXI APB Slave
  // ---------------

  `AXI_ASSIGN(apb_axi_master,master[ariane_soc::APB_SLVS])


  // ---------------
  // AXI hyperbus Slave 
  // ---------------

  axi_cut_intf #(
    .BYPASS     ( 1'b0                     ),
    .ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .USER_WIDTH ( AXI_USER_WIDTH           )
  ) riscvatomics2axihyper_cut (
    .clk_i,
    .rst_ni ( ndmreset_n                ),
    .in     ( hyper_axi_master_cut      ),
    .out    ( hyper_axi_master_redirect )
  );

  `ifdef L3_TCSRAM
  l3_onchip_subsystem # (
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
    ) l3_tcsram (
                                    .clk_i ( clk_i                     ),
                                    .rst_ni( ndmreset_n                ),
                                    .slv   ( hyper_axi_master_redirect )
                                    );
   assign hyper_axi_master.aw_valid = 1'b0;
   assign hyper_axi_master.ar_valid = 1'b0;
   assign hyper_axi_master.w_valid  = 1'b0;
  `else // !`ifdef L3_TCSRAM
    `AXI_ASSIGN(hyper_axi_master,hyper_axi_master_redirect);
  `endif
   
                       
               
  axi_riscv_atomics_wrap #(
    .AXI_ADDR_WIDTH     ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH     ( AXI_DATA_WIDTH           ),
    .AXI_ID_WIDTH       ( ariane_soc::IdWidthSlave ),
    .AXI_USER_WIDTH     ( AXI_USER_WIDTH           ),
    .AXI_MAX_READ_TXNS  ( 8                        ),
    .AXI_MAX_WRITE_TXNS ( 8                        ),
    .RISCV_WORD_WIDTH   ( 64                       )
  ) i_axi_riscv_atomicsl3 (
    .clk_i,
    .rst_ni ( ndmreset_n                ),
    .slv    ( master[ariane_soc::HYAXI] ),
    .mst    ( hyper_axi_master_cut      )
  );
   
  // ---------------
  // AXI CLUSTER Slave
  // ---------------

  `AXI_ASSIGN(cluster_axi_master_cut,master[ariane_soc::Cluster])

  axi_cut_intf #(
    .BYPASS     ( 1'b0                     ),
    .ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .USER_WIDTH ( AXI_USER_WIDTH           )
  ) soc2cluster_cut (
    .clk_i,
    .rst_ni     ( ndmreset_n               ),
    .in         ( cluster_axi_master_cut   ),
    .out        ( cluster_axi_master       )
  );
   
  // ---------------
  // AXI CLUSTER Master
  // ---------------
  `AXI_ASSIGN(slave[ariane_soc::Cluster_Master],cluster_axi_slave)
   
  // ---------------
  // AXI Xbar
  // ---------------
  localparam xbar_cfg_t AXI_XBAR_CFG = '{
                                         NoSlvPorts: ariane_soc::NrSlaves,
                                         NoMstPorts: ariane_soc::NB_PERIPHERALS,
                                         MaxMstTrans: ariane_soc::NB_PERIPHERALS,
                                         MaxSlvTrans: ariane_soc::NrSlaves,
                                         FallThrough: 1'b0,        
                                         LatencyMode: axi_pkg::CUT_ALL_PORTS, // If you cut anything, you might want to remove the soc2cluster_cut.
                                         PipelineStages: 32'd0,
                                         AxiIdWidthSlvPorts: ariane_soc::IdWidth,
                                         AxiIdUsedSlvPorts: ariane_soc::IdWidth,
                                         UniqueIds: 1'b0,
                                         AxiAddrWidth: AXI_ADDRESS_WIDTH,
                                         AxiDataWidth: AXI_DATA_WIDTH,
                                         NoAddrRules: ariane_soc::NB_PERIPHERALS
                                         };

  ariane_soc::addr_map_rule_t [ariane_soc::NB_PERIPHERALS-1:0] addr_map;

 assign addr_map[ariane_soc::Debug] = '{
    idx:  ariane_soc::Debug,
    start_addr: ariane_soc::DebugBase,
    end_addr:   ariane_soc::DebugBase    + ariane_soc::DebugLength  
  };
  assign addr_map[ariane_soc::ROM] = '{ 
    idx:  ariane_soc::ROM,
    start_addr: ariane_soc::ROMBase,
    end_addr:   ariane_soc::ROMBase      + ariane_soc::ROMLength  
  };
  assign addr_map[ariane_soc::UART] = '{ 
    idx:  ariane_soc::UART,
    start_addr: ariane_soc::UARTBase,
    end_addr:   ariane_soc::UARTBase     + ariane_soc::UARTLength  
  };
  assign addr_map[ariane_soc::SERIAL_LINK] = '{ 
    idx:  ariane_soc::SERIAL_LINK,
    start_addr: ariane_soc::SerLink_Base,
    end_addr:   ariane_soc::SerLink_Base + ariane_soc::SerLinkLength  
  };
  assign addr_map[ariane_soc::CLINT] = '{ 
    idx:  ariane_soc::CLINT,
    start_addr: ariane_soc::CLINTBase,
    end_addr:   ariane_soc::CLINTBase    + ariane_soc::CLINTLength  
  };
  assign addr_map[ariane_soc::PLIC] = '{
    idx:  ariane_soc::PLIC,
    start_addr: ariane_soc::PLICBase,
    end_addr:   ariane_soc::PLICBase     + ariane_soc::PLICLength  
  };
  assign addr_map[ariane_soc::Cluster] = '{
    idx:  ariane_soc::Cluster,
    start_addr: ariane_soc::ClusterBase,
    end_addr:   ariane_soc::ClusterBase     + ariane_soc::ClusterLength  
  };
  assign addr_map[ariane_soc::L2SPM] = '{ 
    idx:  ariane_soc::L2SPM,
    start_addr: ariane_soc::L2SPMBase,
    end_addr:   ariane_soc::L2SPMBase     + ariane_soc::L2SPMLength  
  };
  assign addr_map[ariane_soc::APB_SLVS] = '{ 
    idx:  ariane_soc::APB_SLVS,
    start_addr: ariane_soc::APB_SLVSBase,
    end_addr:   ariane_soc::APB_SLVSBase     + ariane_soc::APB_SLVSLength  
  };
  assign addr_map[ariane_soc::Timer] = '{ 
    idx:  ariane_soc::Timer,
    start_addr: ariane_soc::TimerBase,
    end_addr:   ariane_soc::TimerBase    + ariane_soc::TimerLength  
  };
  assign addr_map[ariane_soc::SPI] = '{
    idx:  ariane_soc::SPI,
    start_addr: ariane_soc::SPIBase,
    end_addr:   ariane_soc::SPIBase      + ariane_soc::SPILength  
  };
  assign addr_map[ariane_soc::Ethernet] = '{ 
    idx:  ariane_soc::Ethernet,
    start_addr: ariane_soc::EthernetBase,
    end_addr:   ariane_soc::EthernetBase + ariane_soc::EthernetLength  
  };
  assign addr_map[ariane_soc::HYAXI] = '{ 
    idx:  ariane_soc::HYAXI,
    start_addr: ariane_soc::HYAXIBase,
    end_addr:   ariane_soc::HYAXIBase     + ariane_soc::HYAXILength  
  }; 
  assign addr_map[ariane_soc::AXILiteDom] = '{ 
    idx:  ariane_soc::AXILiteDom,
    start_addr: ariane_soc::AXILiteBase,
    end_addr:   ariane_soc::AXILiteBase + ariane_soc::AXILiteLength  
  }; 

  axi_xbar_intf #(
    .AXI_USER_WIDTH         ( AXI_USER_WIDTH                        ),
    .Cfg                    ( AXI_XBAR_CFG                          ),
    .rule_t                 ( ariane_soc::addr_map_rule_t           )
  ) i_xbar (
    .clk_i                  (clk_i),
    .rst_ni                 (ndmreset_n),
    .test_i                 (1'b0),
    .slv_ports              (slave),
    .mst_ports              (master),
    .addr_map_i             (addr_map),
    .en_default_mst_port_i  ('0), // disable default master port for all slave ports
    .default_mst_port_i     ('0)
  );

  // --------------------
  // AXI Lite Slave    
  // --------------------

  `AXI_ASSIGN(axi_lite_master, master[ariane_soc::AXILiteDom])
   
  // ---------------
  // CLINT
  // ---------------
  // divide clock by two
  logic [3:0] ipi;
  logic [3:0] timer_irq;
  logic rtc_clint;
   
  ariane_axi_soc::req_slv_t    axi_clint_req;
  ariane_axi_soc::resp_slv_t   axi_clint_resp;

  always_ff @(posedge rtc_i or negedge ndmreset_n) begin
    if (~ndmreset_n) begin
      rtc_clint <= 0;
    end else begin
      rtc_clint <= rtc_clint ^ 1'b1;
    end
  end
   
  clint #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH          ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH             ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave   ),
    .lite_req_t     ( ariane_axi_soc::req_slv_t  ),
    .lite_resp_t    ( ariane_axi_soc::resp_slv_t ),
    .NR_CORES       ( 4                          )
  ) i_clint (
    .clk_i       ( clk_i          ),
    .rst_ni      ( ndmreset_n     ),
    .testmode_i  ( test_en        ),
    .axi_req_i   ( axi_clint_req  ),
    .axi_resp_o  ( axi_clint_resp ),
    .rtc_i       ( rtc_clint      ),
    .timer_irq_o ( timer_irq      ),
    .ipi_o       ( ipi            )
  );

  `AXI_ASSIGN_TO_REQ(axi_clint_req,master[ariane_soc::CLINT])
  `AXI_ASSIGN_FROM_RESP(master[ariane_soc::CLINT],axi_clint_resp)


  // ---------------
  // DDR SERIAL LINK
  // ---------------

  ariane_axi_soc::req_t ddr_1_in_req, ddr_1_out_req;
  ariane_axi_soc::resp_t ddr_1_in_rsp, ddr_1_out_rsp;

  logic [3:0] ddr_i, ddr_o;

  localparam RegAw  = 32;
  localparam RegDw  = 32;

  typedef logic [RegAw-1:0]   reg_addr_t;
  typedef logic [RegDw-1:0]   reg_data_t;
  typedef logic [RegDw/8-1:0] reg_strb_t;

  `REG_BUS_TYPEDEF_REQ(reg_req_t, reg_addr_t, reg_data_t, reg_strb_t)
  `REG_BUS_TYPEDEF_RSP(reg_rsp_t, reg_data_t)
 
  reg_req_t   reg_req;
  reg_rsp_t   reg_rsp;

  axi_serializer_intf #(
    .AXI_ID_WIDTH   ( ariane_soc::IdWidthSlave ),
    .MAX_READ_TXNS  ( ariane_soc::NrSlaves     ),
    .MAX_WRITE_TXNS ( ariane_soc::NrSlaves     ),
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH           ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH           )
     )serial_link_serializer (
       .clk_i  ( clk_i                           ),
       .rst_ni ( ndmreset_n                      ),
       .slv    ( master[ariane_soc::SERIAL_LINK] ),
       .mst    ( serial_link_cut                 )
     );

  axi_cut_intf #(
    .BYPASS     ( 1'b0                ),
    .ADDR_WIDTH ( AXI_ADDRESS_WIDTH   ),
    .DATA_WIDTH ( AXI_DATA_WIDTH      ),
    .ID_WIDTH   ( ariane_soc::IdWidth ),
    .USER_WIDTH ( AXI_USER_WIDTH      )
  ) serial_link_cutter (
    .clk_i,
    .rst_ni ( ndmreset_n                ),
    .in     ( serial_link_cut           ),
    .out    ( serial_link_master        )
  );
   
  `AXI_ASSIGN_TO_REQ(ddr_1_in_req,serial_link_master)
  `AXI_ASSIGN_FROM_RESP(serial_link_master, ddr_1_in_rsp)

  `AXI_ASSIGN_FROM_REQ(slave[ariane_soc::Serial_Link], ddr_1_out_req)
  `AXI_ASSIGN_TO_RESP(ddr_1_out_rsp, slave[ariane_soc::Serial_Link])

  `REG_BUS_ASSIGN_TO_REQ(reg_req,serial_linkcfg_reg_master)
  `REG_BUS_ASSIGN_FROM_RSP(serial_linkcfg_reg_master,reg_rsp)

  assign ddr_i[0] = pad_to_serial_link.ddr0_i;
  assign ddr_i[1] = pad_to_serial_link.ddr1_i;
  assign ddr_i[2] = pad_to_serial_link.ddr2_i;
  assign ddr_i[3] = pad_to_serial_link.ddr3_i;

  assign serial_link_to_pad.ddr0_o = ddr_o[0];
  assign serial_link_to_pad.ddr1_o = ddr_o[1];
  assign serial_link_to_pad.ddr2_o = ddr_o[2];
  assign serial_link_to_pad.ddr3_o = ddr_o[3];

   // first serial instance
  serial_link #(
    .axi_req_t        ( ariane_axi_soc::req_t       ),
    .axi_rsp_t        ( ariane_axi_soc::resp_t      ),
    .aw_chan_t        ( ariane_axi_soc::aw_chan_t   ),
    .ar_chan_t        ( ariane_axi_soc::ar_chan_t   ),
    .cfg_req_t        ( reg_req_t   ),
    .cfg_rsp_t        ( reg_rsp_t   )
  ) i_serial_link_1 (
      .clk_i          ( clk_i           ),
      .rst_ni         ( ndmreset_n      ),
      .testmode_i     ( 1'b0            ),
      .axi_in_req_i   ( ddr_1_in_req    ), //slv -> mst axi
      .axi_in_rsp_o   ( ddr_1_in_rsp    ), //slv -> mst axi

      .axi_out_req_o  ( ddr_1_out_req   ), //mst -> slv axi
      .axi_out_rsp_i  ( ddr_1_out_rsp   ), //mst -> slv axi

      .cfg_req_i      ( reg_req ), //reg_req from apb slave
      .cfg_rsp_o      ( reg_rsp ), //reg_rsp apb slave
      
      .ddr_clk_i      ( pad_to_serial_link.ddr_clk_i ),
      .ddr_i          ( ddr_i ),
      .ddr_o          ( ddr_o )
  );



  // ---------------
  // Peripherals
  // ---------------
  logic tx, rx;
  logic [7:0] irqs;

  ariane_peripherals #(
    .AxiAddrWidth ( AXI_ADDRESS_WIDTH        ),
    .AxiDataWidth ( AXI_DATA_WIDTH           ),
    .AxiIdWidth   ( ariane_soc::IdWidthSlave ),
`ifdef PMU_BLOCK
    .PMU_NUM_COUNTER  ( PMU_NUM_COUNTER      ),
`endif    
`ifdef TARGET_SYNTHESIS
    .InclUART     ( 1'b1                     ),
`else
    .InclUART     ( 1'b0                     ),
`endif
`ifdef TARGET_FPGA  
    .InclSPI      ( 1'b1                     ),
`else
    .InclSPI      ( 1'b0                     ),
`endif
    .InclEthernet ( 1'b0                     )
  ) i_ariane_peripherals (
    .clk_i           ( clk_i                        ),
    .rst_ni          ( ndmreset_n                   ),
    .plic            ( master[ariane_soc::PLIC]     ),
    .uart            ( master[ariane_soc::UART]     ),
    .spi             ( master[ariane_soc::SPI]      ),
    .ethernet        ( master[ariane_soc::Ethernet] ),
    .timer           ( master[ariane_soc::Timer]    ),
    .udma_evt_i      ( udma_events_i                ),
    .cluster_eoc_i   ( cluster_eoc_i                ),
    .c2h_irq_i       ( c2h_irq_i                    ),
    .can_irq_i       ( can_irq_i                    ),
    .cl_dma_pe_evt_i ( cl_dma_pe_evt_i              ),
    .irq_o           ( irqs                         ),
    .rx_i            ( cva6_uart_rx_i               ),
    .tx_o            ( cva6_uart_tx_o               ),

    `ifdef PMU_BLOCK
    .pmu_intr_i      ( pmu_intr_i                   ),
    `endif

    .eth_txck        ( ),
    .eth_rxck        ( ),
    .eth_rxctl       ( ),
    .eth_rxd         ( ),
    .eth_rst_n       ( ),
    .eth_tx_en       ( ),
    .eth_txd         ( ),
    .phy_mdio        ( ),
    .eth_mdc         ( ),
    .mdio            ( ),
    .mdc             ( )
  );

  // --------------------
  // SPUs on cores output
  // --------------------

  localparam N_ADDR_RULES = 2;
  ariane_soc::addr_map_rule_t [N_ADDR_RULES-1:0]   spu_core_addr_map;
  assign spu_core_addr_map[0] = '{
        idx: 0,
        start_addr: ariane_soc::DebugBase,
        end_addr:   ariane_soc::HYAXIBase
  };

  assign spu_core_addr_map[1] = '{
        idx: 1,
        start_addr: ariane_soc::HYAXIBase,
        end_addr:   ariane_soc::HYAXIBase + ariane_soc::HYAXILength
  };

  spu_top #(
    // Static configuration parameters of the cache.
    .SetAssociativity   ( ariane_soc::LLC_SET_ASSOC   ),
    .NumLines           ( ariane_soc::LLC_NUM_LINES   ),
    .NumBlocks          ( ariane_soc::LLC_NUM_BLOCKS  ),
    // AXI4 Specifications
    .IdWidthMasters     ( ariane_soc::IdWidth         ),
    .IdWidthSlaves      ( ariane_soc::IdWidthSlave+ 1 ),
    .AddrWidth          ( AXI_ADDRESS_WIDTH           ),
    .DataWidth          ( AXI_DATA_WIDTH              ),
    // Address Indexing
    .addr_rule_t        ( ariane_soc::addr_map_rule_t ),
    .N_ADDR_RULES       ( N_ADDR_RULES                ),
    // FIFO and CAM Parameters
    .CAM_DEPTH          (  3                          ),
    .FIFO_DEPTH         (  3                          )
  ) i_spu_core_0_llc (
    .clk_i              ( clk_i                       ),
    .rst_ni             ( rst_ni                      ),
    .addr_map_i         ( spu_core_addr_map           ),
    .spu_slv            ( slave_to_spu[ariane_soc::Core_0-4] ),
    .spu_mst            ( slave[ariane_soc::Core_0]   ),
    .e_out              ( spu_core_0_out              )
  );

  spu_top #(
    // Static configuration parameters of the cache.
    .SetAssociativity   ( ariane_soc::LLC_SET_ASSOC   ),
    .NumLines           ( ariane_soc::LLC_NUM_LINES   ),
    .NumBlocks          ( ariane_soc::LLC_NUM_BLOCKS  ),
    // AXI4 Specifications
    .IdWidthMasters     ( ariane_soc::IdWidth         ),
    .IdWidthSlaves      ( ariane_soc::IdWidthSlave+ 1 ),
    .AddrWidth          ( AXI_ADDRESS_WIDTH           ),
    .DataWidth          ( AXI_DATA_WIDTH              ),
    // Address Indexing
    .addr_rule_t        ( ariane_soc::addr_map_rule_t ),
    .N_ADDR_RULES       ( N_ADDR_RULES                ),
    // FIFO and CAM Parameters
    .CAM_DEPTH          (  3                          ),
    .FIFO_DEPTH         (  3                          )
  ) i_spu_core_1_llc (
    .clk_i              ( clk_i                       ),
    .rst_ni             ( rst_ni                      ),
    .addr_map_i         ( spu_core_addr_map           ),
    .spu_slv            ( slave_to_spu[ariane_soc::Core_1-4] ),
    .spu_mst            ( slave[ariane_soc::Core_1]   ),
    .e_out              ( spu_core_1_out              )
  );

  spu_top #(
    // Static configuration parameters of the cache.
    .SetAssociativity   ( ariane_soc::LLC_SET_ASSOC   ),
    .NumLines           ( ariane_soc::LLC_NUM_LINES   ),
    .NumBlocks          ( ariane_soc::LLC_NUM_BLOCKS  ),
    // AXI4 Specifications
    .IdWidthMasters     ( ariane_soc::IdWidth         ),
    .IdWidthSlaves      ( ariane_soc::IdWidthSlave+ 1 ),
    .AddrWidth          ( AXI_ADDRESS_WIDTH           ),
    .DataWidth          ( AXI_DATA_WIDTH              ),
    // Address Indexing
    .addr_rule_t        ( ariane_soc::addr_map_rule_t ),
    .N_ADDR_RULES       ( N_ADDR_RULES                ),
    // FIFO and CAM Parameters
    .CAM_DEPTH          (  3                          ),
    .FIFO_DEPTH         (  3                          )
  ) i_spu_core_2_llc (
    .clk_i              ( clk_i                       ),
    .rst_ni             ( rst_ni                      ),
    .addr_map_i         ( spu_core_addr_map           ),
    .spu_slv            ( slave_to_spu[ariane_soc::Core_2-4] ),
    .spu_mst            ( slave[ariane_soc::Core_2]   ),
    .e_out              ( spu_core_2_out              )
  );

  spu_top #(
    // Static configuration parameters of the cache.
    .SetAssociativity   ( ariane_soc::LLC_SET_ASSOC   ),
    .NumLines           ( ariane_soc::LLC_NUM_LINES   ),
    .NumBlocks          ( ariane_soc::LLC_NUM_BLOCKS  ),
    // AXI4 Specifications
    .IdWidthMasters     ( ariane_soc::IdWidth         ),
    .IdWidthSlaves      ( ariane_soc::IdWidthSlave+ 1 ),
    .AddrWidth          ( AXI_ADDRESS_WIDTH           ),
    .DataWidth          ( AXI_DATA_WIDTH              ),
    // Address Indexing
    .addr_rule_t        ( ariane_soc::addr_map_rule_t ),
    .N_ADDR_RULES       ( N_ADDR_RULES                ),
    // FIFO and CAM Parameters
    .CAM_DEPTH          (  3                          ),
    .FIFO_DEPTH         (  3                          )
  ) i_spu_core_3_llc (
    .clk_i              ( clk_i                       ),
    .rst_ni             ( rst_ni                      ),
    .addr_map_i         ( spu_core_addr_map           ),
    .spu_slv            ( slave_to_spu[ariane_soc::Core_3-4] ),
    .spu_mst            ( slave[ariane_soc::Core_3]   ),
    .e_out              ( spu_core_3_out              )
  );
  // ---------------
  // Core #0
  // ---------------

  cva6_synth_wrap #(
    .LOG_DEPTH (1)
  ) i_ariane_wrap_0 (
    .clk_i                ( cva6_clk_i                    ),
    .rst_ni               ( cva6_rst_ni                   ),
    .boot_addr_i          ( ariane_soc::ROMBase           ), // start fetching from ROM
    .hart_id_i            ( 64'd0                         ),
    .irq_i                ( irqs[1:0]                     ), // async signal
    .ipi_i                ( ipi[0]                        ), // async signal
    .time_irq_i           ( timer_irq[0]                  ), // async signal
    .debug_req_i          ( debug_req_core[0]             ), // async signal
    .data_master_aw_wptr_o( cva6_axi_master_dst_0.aw_wptr ),
    .data_master_aw_data_o( cva6_axi_master_dst_0.aw_data ), 
    .data_master_aw_rptr_i( cva6_axi_master_dst_0.aw_rptr ),
    .data_master_ar_wptr_o( cva6_axi_master_dst_0.ar_wptr ),
    .data_master_ar_data_o( cva6_axi_master_dst_0.ar_data ),
    .data_master_ar_rptr_i( cva6_axi_master_dst_0.ar_rptr ),
    .data_master_w_wptr_o ( cva6_axi_master_dst_0.w_wptr  ),
    .data_master_w_data_o ( cva6_axi_master_dst_0.w_data  ),
    .data_master_w_rptr_i ( cva6_axi_master_dst_0.w_rptr  ),
    .data_master_r_wptr_i ( cva6_axi_master_dst_0.r_wptr  ),
    .data_master_r_data_i ( cva6_axi_master_dst_0.r_data  ),
    .data_master_r_rptr_o ( cva6_axi_master_dst_0.r_rptr  ),
    .data_master_b_wptr_i ( cva6_axi_master_dst_0.b_wptr  ),
    .data_master_b_data_i ( cva6_axi_master_dst_0.b_data  ),
    .data_master_b_rptr_o ( cva6_axi_master_dst_0.b_rptr  )
  );

  axi_cdc_dst_intf #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH         ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH            ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth       ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH            ),
    .LOG_DEPTH      ( 1                         )
  ) cva6_0_to_xbar (
    .src            ( cva6_axi_master_dst_0     ),
    .dst_clk_i      ( clk_i                     ),
    .dst_rst_ni     ( ndmreset_n                ),
  `ifdef PMU_BLOCK
    .dst            ( slave_to_spu[ariane_soc::Core_0-4] )
  `else
    .dst            ( slave[ariane_soc::Core_0] )
  `endif
  );

  // ---------------
  // Core #1
  // ---------------

  cva6_synth_wrap #(
    .LOG_DEPTH (1)
  ) i_ariane_wrap_1 (
    .clk_i                ( cva6_clk_i                    ),
    .rst_ni               ( cva6_rst_ni                   ),
    .boot_addr_i          ( ariane_soc::ROMBase           ), // start fetching from ROM
    .hart_id_i            ( 64'd1                         ),
    .irq_i                ( irqs[3:2]                     ), // async signal
    .ipi_i                ( ipi[1]                        ), // async signal
    .time_irq_i           ( timer_irq[1]                  ), // async signal
    .debug_req_i          ( debug_req_core[1]             ), // async signal
    .data_master_aw_wptr_o( cva6_axi_master_dst_1.aw_wptr ),
    .data_master_aw_data_o( cva6_axi_master_dst_1.aw_data ), 
    .data_master_aw_rptr_i( cva6_axi_master_dst_1.aw_rptr ),
    .data_master_ar_wptr_o( cva6_axi_master_dst_1.ar_wptr ),
    .data_master_ar_data_o( cva6_axi_master_dst_1.ar_data ),
    .data_master_ar_rptr_i( cva6_axi_master_dst_1.ar_rptr ),
    .data_master_w_wptr_o ( cva6_axi_master_dst_1.w_wptr  ),
    .data_master_w_data_o ( cva6_axi_master_dst_1.w_data  ),
    .data_master_w_rptr_i ( cva6_axi_master_dst_1.w_rptr  ),
    .data_master_r_wptr_i ( cva6_axi_master_dst_1.r_wptr  ),
    .data_master_r_data_i ( cva6_axi_master_dst_1.r_data  ),
    .data_master_r_rptr_o ( cva6_axi_master_dst_1.r_rptr  ),
    .data_master_b_wptr_i ( cva6_axi_master_dst_1.b_wptr  ),
    .data_master_b_data_i ( cva6_axi_master_dst_1.b_data  ),
    .data_master_b_rptr_o ( cva6_axi_master_dst_1.b_rptr  )
  );

  axi_cdc_dst_intf #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH         ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH            ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth       ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH            ),
    .LOG_DEPTH      ( 1                         )
  ) cva6_1_to_xbar (
    .src            ( cva6_axi_master_dst_1     ),
    .dst_clk_i      ( clk_i                     ),
    .dst_rst_ni     ( ndmreset_n                ),
  `ifdef PMU_BLOCK
    .dst            ( slave_to_spu[ariane_soc::Core_1-4] )
  `else
    .dst            ( slave[ariane_soc::Core_1] )
  `endif
  );

  // ---------------
  // Core #2
  // ---------------

  cva6_synth_wrap #(
    .LOG_DEPTH (1)
  ) i_ariane_wrap_2 (
    .clk_i                ( cva6_clk_i                    ),
    .rst_ni               ( cva6_rst_ni                   ),
    .boot_addr_i          ( ariane_soc::ROMBase           ), // start fetching from ROM
    .hart_id_i            ( 64'd2                         ),
    .irq_i                ( irqs[5:4]                     ), // async signal
    .ipi_i                ( ipi[2]                        ), // async signal
    .time_irq_i           ( timer_irq[2]                  ), // async signal
    .debug_req_i          ( debug_req_core[2]             ), // async signal
    .data_master_aw_wptr_o( cva6_axi_master_dst_2.aw_wptr ),
    .data_master_aw_data_o( cva6_axi_master_dst_2.aw_data ), 
    .data_master_aw_rptr_i( cva6_axi_master_dst_2.aw_rptr ),
    .data_master_ar_wptr_o( cva6_axi_master_dst_2.ar_wptr ),
    .data_master_ar_data_o( cva6_axi_master_dst_2.ar_data ),
    .data_master_ar_rptr_i( cva6_axi_master_dst_2.ar_rptr ),
    .data_master_w_wptr_o ( cva6_axi_master_dst_2.w_wptr  ),
    .data_master_w_data_o ( cva6_axi_master_dst_2.w_data  ),
    .data_master_w_rptr_i ( cva6_axi_master_dst_2.w_rptr  ),
    .data_master_r_wptr_i ( cva6_axi_master_dst_2.r_wptr  ),
    .data_master_r_data_i ( cva6_axi_master_dst_2.r_data  ),
    .data_master_r_rptr_o ( cva6_axi_master_dst_2.r_rptr  ),
    .data_master_b_wptr_i ( cva6_axi_master_dst_2.b_wptr  ),
    .data_master_b_data_i ( cva6_axi_master_dst_2.b_data  ),
    .data_master_b_rptr_o ( cva6_axi_master_dst_2.b_rptr  )
  );

  axi_cdc_dst_intf #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH         ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH            ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth       ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH            ),
    .LOG_DEPTH      ( 1                         )
  ) cva6_2_to_xbar (
    .src            ( cva6_axi_master_dst_2     ),
    .dst_clk_i      ( clk_i                     ),
    .dst_rst_ni     ( ndmreset_n                ),
  `ifdef PMU_BLOCK
    .dst            ( slave_to_spu[ariane_soc::Core_2-4] )
  `else
    .dst            ( slave[ariane_soc::Core_2] )
  `endif
  );

  // // ---------------
  // // Core #3
  // // ---------------

  cva6_synth_wrap #(
    .LOG_DEPTH (1)
  ) i_ariane_wrap_3 (
    .clk_i                ( cva6_clk_i                    ),
    .rst_ni               ( cva6_rst_ni                   ),
    .boot_addr_i          ( ariane_soc::ROMBase           ), // start fetching from ROM
    .hart_id_i            ( 64'd3                         ),
    .irq_i                ( irqs[7:6]                     ), // async signal
    .ipi_i                ( ipi[3]                        ), // async signal
    .time_irq_i           ( timer_irq[3]                  ), // async signal
    .debug_req_i          ( debug_req_core[3]             ), // async signal
    .data_master_aw_wptr_o( cva6_axi_master_dst_3.aw_wptr ),
    .data_master_aw_data_o( cva6_axi_master_dst_3.aw_data ), 
    .data_master_aw_rptr_i( cva6_axi_master_dst_3.aw_rptr ),
    .data_master_ar_wptr_o( cva6_axi_master_dst_3.ar_wptr ),
    .data_master_ar_data_o( cva6_axi_master_dst_3.ar_data ),
    .data_master_ar_rptr_i( cva6_axi_master_dst_3.ar_rptr ),
    .data_master_w_wptr_o ( cva6_axi_master_dst_3.w_wptr  ),
    .data_master_w_data_o ( cva6_axi_master_dst_3.w_data  ),
    .data_master_w_rptr_i ( cva6_axi_master_dst_3.w_rptr  ),
    .data_master_r_wptr_i ( cva6_axi_master_dst_3.r_wptr  ),
    .data_master_r_data_i ( cva6_axi_master_dst_3.r_data  ),
    .data_master_r_rptr_o ( cva6_axi_master_dst_3.r_rptr  ),
    .data_master_b_wptr_i ( cva6_axi_master_dst_3.b_wptr  ),
    .data_master_b_data_i ( cva6_axi_master_dst_3.b_data  ),
    .data_master_b_rptr_o ( cva6_axi_master_dst_3.b_rptr  )
  );

  axi_cdc_dst_intf #(
    .AXI_ADDR_WIDTH ( AXI_ADDRESS_WIDTH         ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH            ),
    .AXI_ID_WIDTH   ( ariane_soc::IdWidth       ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH            ),
    .LOG_DEPTH      ( 1                         )
  ) cva6_3_to_xbar (
    .src            ( cva6_axi_master_dst_3     ),
    .dst_clk_i      ( clk_i                     ),
    .dst_rst_ni     ( ndmreset_n                ),
  `ifdef PMU_BLOCK
    .dst            ( slave_to_spu[ariane_soc::Core_3-4] )
  `else
    .dst            ( slave[ariane_soc::Core_3] )
  `endif
  );
   
endmodule
